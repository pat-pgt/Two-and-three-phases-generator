library IEEE;
use IEEE.Std_Logic_1164.all,
ieee.numeric_std.all,
work.cmos74hc.all;

package super_triphase is
  component super_triphase_gene is
    port(
      signal CLK : in std_logic;
      SIGNAL P4_Q7 : out Std_Logic;
      SIGNAL P4_Q6 : out Std_Logic;
      SIGNAL P4_Q5 : out Std_Logic;
      SIGNAL P4_Q4 : out Std_Logic;
      SIGNAL P4_Q3 : out Std_Logic;
      SIGNAL P4_Q2 : out Std_Logic;
      SIGNAL P4_Q1 : out Std_Logic;
      SIGNAL P4_Q0 : out Std_Logic;
      SIGNAL P1_Q7 : out Std_Logic;
      SIGNAL P1_Q6 : out Std_Logic;
      SIGNAL P1_Q5 : out Std_Logic;
      SIGNAL P1_Q4 : out Std_Logic;
      SIGNAL P1_Q3 : out Std_Logic;
      SIGNAL P1_Q2 : out Std_Logic;
      SIGNAL P1_Q1 : out Std_Logic;
      SIGNAL P1_Q0 : out Std_Logic;
      SIGNAL P2_Q7 : out Std_Logic;
      SIGNAL P2_Q6 : out Std_Logic;
      SIGNAL P2_Q5 : out Std_Logic;
      SIGNAL P2_Q4 : out Std_Logic;
      SIGNAL P2_Q3 : out Std_Logic;
      SIGNAL P2_Q2 : out Std_Logic;
      SIGNAL P2_Q1 : out Std_Logic;
      SIGNAL P2_Q0 : out Std_Logic;
      SIGNAL P3_Q7 : out Std_Logic;
      SIGNAL P3_Q6 : out Std_Logic;
      SIGNAL P3_Q5 : out Std_Logic;
      SIGNAL P3_Q4 : out Std_Logic;
      SIGNAL P3_Q3 : out Std_Logic;
      SIGNAL P3_Q2 : out Std_Logic;
      SIGNAL P3_Q1 : out Std_Logic;
      SIGNAL P3_Q0 : out Std_Logic);
  end component super_triphase_gene;
end package super_triphase;

-- Structural VHDL generated by gnetlist
-- Context clause
library IEEE;
use IEEE.Std_Logic_1164.all,
  ieee.numeric_std.all,
  work.cmos74hc.all;
-- Entity declaration

ENTITY super_triphase_gene IS
  port (
    signal CLK : in std_logic;
    SIGNAL P4_Q7 : out Std_Logic;
    SIGNAL P4_Q6 : out Std_Logic;
    SIGNAL P4_Q5 : out Std_Logic;
    SIGNAL P4_Q4 : out Std_Logic;
    SIGNAL P4_Q3 : out Std_Logic;
    SIGNAL P4_Q2 : out Std_Logic;
    SIGNAL P4_Q1 : out Std_Logic;
      SIGNAL P4_Q0 : out Std_Logic;
      SIGNAL P1_Q7 : out Std_Logic;
      SIGNAL P1_Q6 : out Std_Logic;
      SIGNAL P1_Q5 : out Std_Logic;
      SIGNAL P1_Q4 : out Std_Logic;
      SIGNAL P1_Q3 : out Std_Logic;
      SIGNAL P1_Q2 : out Std_Logic;
      SIGNAL P1_Q1 : out Std_Logic;
      SIGNAL P1_Q0 : out Std_Logic;
      SIGNAL P2_Q7 : out Std_Logic;
      SIGNAL P2_Q6 : out Std_Logic;
      SIGNAL P2_Q5 : out Std_Logic;
      SIGNAL P2_Q4 : out Std_Logic;
      SIGNAL P2_Q3 : out Std_Logic;
      SIGNAL P2_Q2 : out Std_Logic;
      SIGNAL P2_Q1 : out Std_Logic;
      SIGNAL P2_Q0 : out Std_Logic;
      SIGNAL P3_Q7 : out Std_Logic;
      SIGNAL P3_Q6 : out Std_Logic;
      SIGNAL P3_Q5 : out Std_Logic;
      SIGNAL P3_Q4 : out Std_Logic;
      SIGNAL P3_Q3 : out Std_Logic;
      SIGNAL P3_Q2 : out Std_Logic;
      SIGNAL P3_Q1 : out Std_Logic;
      SIGNAL P3_Q0 : out Std_Logic);
END super_triphase_gene;


-- Secondary unit
ARCHITECTURE netlist OF super_triphase_gene IS
  
  SIGNAL unnamed_net90 : Std_Logic;
  SIGNAL unnamed_net89 : Std_Logic;
  SIGNAL unnamed_net88 : Std_Logic;
  SIGNAL unnamed_net87 : Std_Logic;
  SIGNAL unnamed_net86 : Std_Logic;
  SIGNAL unnamed_net85 : Std_Logic;
  SIGNAL unnamed_net84 : Std_Logic;
  SIGNAL unnamed_net83 : Std_Logic;
  SIGNAL unnamed_net82 : Std_Logic;
  SIGNAL unnamed_net81 : Std_Logic;
  SIGNAL unnamed_net80 : Std_Logic;
  SIGNAL unnamed_net79 : Std_Logic;
  SIGNAL unnamed_net78 : Std_Logic;
  SIGNAL unnamed_net77 : Std_Logic;
  SIGNAL unnamed_net76 : Std_Logic;
  SIGNAL unnamed_net75 : Std_Logic;
  SIGNAL unnamed_net74 : Std_Logic;
  SIGNAL unnamed_net73 : Std_Logic;
  SIGNAL unnamed_net72 : Std_Logic;
  SIGNAL unnamed_net71 : Std_Logic;
  SIGNAL unnamed_net70 : Std_Logic;
  SIGNAL unnamed_net69 : Std_Logic;
  SIGNAL unnamed_net68 : Std_Logic;
  SIGNAL unnamed_net67 : Std_Logic;
  SIGNAL unnamed_net66 : Std_Logic;
  SIGNAL unnamed_net65 : Std_Logic;
  SIGNAL unnamed_net64 : Std_Logic;
  SIGNAL unnamed_net63 : Std_Logic;
  SIGNAL unnamed_net62 : Std_Logic;
  SIGNAL unnamed_net61 : Std_Logic;
  SIGNAL unnamed_net60 : Std_Logic;
  SIGNAL unnamed_net59 : Std_Logic;
  SIGNAL unnamed_net58 : Std_Logic;
  SIGNAL unnamed_net57 : Std_Logic;
  SIGNAL unnamed_net56 : Std_Logic;
  SIGNAL unnamed_net55 : Std_Logic;
  SIGNAL unnamed_net54 : Std_Logic;
  SIGNAL unnamed_net53 : Std_Logic;
  SIGNAL unnamed_net52 : Std_Logic;
  SIGNAL unnamed_net51 : Std_Logic;
  SIGNAL unnamed_net50 : Std_Logic;
  SIGNAL unnamed_net49 : Std_Logic;
  SIGNAL unnamed_net48 : Std_Logic;

  SIGNAL unnamed_net47 : Std_Logic;
  SIGNAL unnamed_net46 : Std_Logic;
  SIGNAL unnamed_net45 : Std_Logic;
  
  SIGNAL unnamed_net44 : Std_Logic;
  
  SIGNAL unnamed_net43 : Std_Logic;
  
  SIGNAL unnamed_net42 : Std_Logic;
  
  SIGNAL unnamed_net41 : Std_Logic;
  SIGNAL unnamed_net40 : Std_Logic;
  SIGNAL unnamed_net39 : Std_Logic;
  SIGNAL unnamed_net38 : Std_Logic;
  SIGNAL unnamed_net37 : Std_Logic;
  SIGNAL unnamed_net36 : Std_Logic;
  SIGNAL unnamed_net35 : Std_Logic;
  SIGNAL unnamed_net34 : Std_Logic;
  SIGNAL unnamed_net33 : Std_Logic;
  SIGNAL unnamed_net32 : Std_Logic;
  SIGNAL unnamed_net31 : Std_Logic;
  SIGNAL unnamed_net30 : Std_Logic;
  SIGNAL unnamed_net29 : Std_Logic;
  SIGNAL unnamed_net28 : Std_Logic;
  SIGNAL unnamed_net27 : Std_Logic;
  SIGNAL unnamed_net26 : Std_Logic;
  SIGNAL unnamed_net25 : Std_Logic;
  SIGNAL unnamed_net24 : Std_Logic;
  SIGNAL unnamed_net23 : Std_Logic;
  SIGNAL unnamed_net22 : Std_Logic;
  SIGNAL unnamed_net21 : Std_Logic;
  SIGNAL unnamed_net20 : Std_Logic;
  SIGNAL unnamed_net19 : Std_Logic;
  SIGNAL unnamed_net18 : Std_Logic;
  SIGNAL unnamed_net17 : Std_Logic;
  SIGNAL unnamed_net16 : Std_Logic;
  SIGNAL unnamed_net15 : Std_Logic;
  SIGNAL unnamed_net14 : Std_Logic;
  SIGNAL unnamed_net13 : Std_Logic;
  SIGNAL unnamed_net12 : Std_Logic;
  SIGNAL unnamed_net11 : Std_Logic;
  SIGNAL Vcc : Std_Logic;
  SIGNAL GND : Std_Logic;
  SIGNAL unnamed_net10 : Std_Logic;
  SIGNAL unnamed_net9 : Std_Logic;
  SIGNAL unnamed_net8 : Std_Logic;
  SIGNAL unnamed_net7 : Std_Logic;
  SIGNAL unnamed_net6 : Std_Logic;
  SIGNAL unnamed_net5 : Std_Logic;
  SIGNAL unnamed_net4 : Std_Logic;
  SIGNAL unnamed_net3 : Std_Logic;
  SIGNAL unnamed_net2 : Std_Logic;
  SIGNAL unnamed_net1 : Std_Logic;
BEGIN
-- Architecture statement part
  U23 : hc7485
    PORT MAP (
      P10 => unnamed_net79,
      P5 => unnamed_net88,
      P12 => unnamed_net80,
      P6 => unnamed_net89,
      P13 => GND,
      P7 => unnamed_net90,
      P15 => GND,
      P9 => unnamed_net28,
      P11 => unnamed_net29,
      P14 => GND,
      P1 => GND,
      P4 => GND,
      P3 => GND,
      P2 => GND,
      P16 => Vcc,
      P8 => GND);

  U22 : hc7485
    PORT MAP (
      P10 => unnamed_net81,
      P5 => unnamed_net86,
      P12 => unnamed_net83,
      P6 => unnamed_net87,
      P13 => unnamed_net82,
      P7 => unnamed_net47,
      P15 => unnamed_net78,
      P9 => unnamed_net30,
      P11 => unnamed_net31,
      P14 => unnamed_net32,
      P1 => unnamed_net33,
      P4 => unnamed_net88,
      P3 => unnamed_net89,
      P2 => unnamed_net90,
      P16 => Vcc,
      P8 => GND);

  U21 : hc7420
    PORT MAP (
      P6 => unnamed_net81,
      P5 => unnamed_net73,
      P1 => unnamed_net68,
      P2 => unnamed_net72,
      P4 => unnamed_net73,
      
      P8 => unnamed_net83,
      P13 => unnamed_net75,
      P9 => unnamed_net72,
      P10 => unnamed_net70,
      P12 => unnamed_net74,
      P14 => Vcc,
      P7 => GND);

  U20 : hc7400
    PORT MAP (
      P3 => unnamed_net78,
      P2 => unnamed_net75,
      P1 => unnamed_net58,
      
      P6 => unnamed_net79,
      P5 => unnamed_net73,
      P4 => unnamed_net67,
      
      P8 => unnamed_net80,
      P10 => unnamed_net81,
      P9 => unnamed_net72,
      
      P11 => unnamed_net82,
      P13 => unnamed_net74,
      P12 => unnamed_net73,
      P14 => Vcc,
      P7 => GND);

  U18 : hc74163
    PORT MAP (
      P3 => GND,
      P14 => unnamed_net67,
      P4 => GND,
      P13 => unnamed_net69,
      P5 => GND,
      P12 => unnamed_net71,
      P6 => GND,
      P11 => unnamed_net76,
      P7 => Vcc,
      P15 => unnamed_net77,
      P10 => Vcc,
      P2 => CLK,
      P1 => Vcc,
      P9 => unnamed_net48,
      P16 => Vcc,
      P8 => GND);

  U19 : hc74138
    PORT MAP (
      P1 => unnamed_net67,
      P15 => unnamed_net68,
      P2 => unnamed_net69,
      P14 => unnamed_net70,
      P3 => unnamed_net71,
      P13 => unnamed_net72,
      P12 => unnamed_net73,
      P4 => GND,
      P11 => unnamed_net74,
      P5 => GND,
      P10 => unnamed_net58,
      P6 => Vcc,
      P9 => unnamed_net75,
      P7 => unnamed_net48,
      P16 => Vcc,
      P8 => GND);

  U17 : hc7473
    PORT MAP (
      P14 => unnamed_net57,
      P12 => unnamed_net27,
      P3 => unnamed_net58,
      P13 => unnamed_net65,
      P2 => Vcc,
      P1 => CLK,
      
      P7 => GND,
      P9 => unnamed_net84,
      P10 => GND,
      P8 => unnamed_net85,
      P6 => GND,
      P5 => GND,
      P4 => Vcc,
      P11 => GND);

  U16 : hc7473
    PORT MAP (
      P14 => unnamed_net27,
      P12 => unnamed_net64,
      P3 => unnamed_net65,
      P13 => unnamed_net60,
      P2 => Vcc,
      P1 => CLK,
      
      P7 => unnamed_net64,
      P9 => unnamed_net66,
      P10 => unnamed_net60,
      P8 => unnamed_net21,
      P6 => Vcc,
      P5 => CLK,
      P4 => Vcc,
      P11 => GND);

  U8 : hc74138
    PORT MAP (
      P1 => unnamed_net22,
      P15 => unnamed_net42,
      P2 => unnamed_net23,
      P14 => unnamed_net43,
      P3 => GND,
      P13 => unnamed_net40,
      P12 => unnamed_net44,
      P4 => GND,
      P11 => unnamed_net59,
      P5 => unnamed_net60,
      P10 => unnamed_net61,
      P6 => Vcc,
      P9 => unnamed_net62,
      P7 => unnamed_net63,
      P16 => Vcc,
      P8 => GND);

  U7 : hc7400
    PORT MAP (
      P8 => unnamed_net9,
      P10 => unnamed_net55,
      P9 => unnamed_net56,
      
      P11 => unnamed_net56,
      P13 => unnamed_net23,
      P12 => Vcc,
      
      P3 => unnamed_net20,
      P2 => unnamed_net56,
      P1 => unnamed_net22,
      
      P6 => unnamed_net57,
      P5 => Vcc,
      P4 => unnamed_net58,
      P14 => Vcc,
      P7 => GND);

  U3 : hc74163
    PORT MAP (
      P3 => GND,
      P14 => unnamed_net49,
      P4 => Vcc,
      P13 => unnamed_net50,
      P5 => GND,
      P12 => unnamed_net51,
      P6 => Vcc,
      P11 => unnamed_net52,
      P7 => Vcc,
      P15 => unnamed_net53,
      P10 => Vcc,
      P2 => CLK,
      P1 => Vcc,
      P9 => unnamed_net54,
      P16 => Vcc,
      P8 => GND);

  U2 : hc74163
    PORT MAP (
      P3 => GND,
      P14 => unnamed_net38,
      P4 => GND,
      P13 => unnamed_net36,
      P5 => GND,
      P12 => unnamed_net34,
      P6 => GND,
      P11 => unnamed_net45,
      P7 => Vcc,
      P15 => unnamed_net46,
      P10 => unnamed_net47,
      P2 => CLK,
      P1 => Vcc,
      P9 => unnamed_net48,
      P16 => Vcc,
      P8 => GND);

  U15 : hc74273
    PORT MAP (
      P11 => unnamed_net44,
      P3 => unnamed_net39,
      P4 => unnamed_net37,
      P7 => unnamed_net35,
      P8 => unnamed_net35,
      P13 => unnamed_net41,
      P14 => unnamed_net41,
      P17 => unnamed_net41,
      P18 => unnamed_net41,
      P1 => Vcc,
      P2 => P4_Q0,
      P5 => P4_Q1,
      P6 => P4_Q2,
      P9 => P4_Q3,
      P12 => P4_Q4,
      P15 => P4_Q5,
      P16 => P4_Q6,
      P19 => P4_Q7,
      P20 => Vcc,
      P10 => GND);

  U12 : hc74273
    PORT MAP (
      P11 => unnamed_net43,
      P3 => unnamed_net39,
      P4 => unnamed_net37,
      P7 => unnamed_net35,
      P8 => unnamed_net35,
      P13 => unnamed_net41,
      P14 => unnamed_net41,
      P17 => unnamed_net41,
      P18 => unnamed_net41,
      P1 => Vcc,
      P2 => P1_Q0,
      P5 => P1_Q1,
      P6 => P1_Q2,
      P9 => P1_Q3,
      P12 => P1_Q4,
      P15 => P1_Q5,
      P16 => P1_Q6,
      P19 => P1_Q7,
      P20 => Vcc,
      P10 => GND);

  U13 : hc74273
    PORT MAP (
      P11 => unnamed_net42,
      P3 => unnamed_net39,
      P4 => unnamed_net37,
      P7 => unnamed_net35,
      P8 => unnamed_net35,
      P13 => unnamed_net41,
      P14 => unnamed_net41,
      P17 => unnamed_net41,
      P18 => unnamed_net41,
      P1 => Vcc,
      P2 => P2_Q0,
      P5 => P2_Q1,
      P6 => P2_Q2,
      P9 => P2_Q3,
      P12 => P2_Q4,
      P15 => P2_Q5,
      P16 => P2_Q6,
      P19 => P2_Q7,
      P20 => Vcc,
      P10 => GND);

  U14 : hc74273
    PORT MAP (
      P11 => unnamed_net40,
      P3 => unnamed_net39,
      P4 => unnamed_net37,
      P7 => unnamed_net35,
      P8 => unnamed_net35,
      P13 => unnamed_net41,
      P14 => unnamed_net41,
      P17 => unnamed_net41,
      P18 => unnamed_net41,
      P1 => Vcc,
      P2 => P3_Q0,
      P5 => P3_Q1,
      P6 => P3_Q2,
      P9 => P3_Q3,
      P12 => P3_Q4,
      P15 => P3_Q5,
      P16 => P3_Q6,
      P19 => P3_Q7,
      P20 => Vcc,
      P10 => GND);

  U11 : hc7486
    PORT MAP (
      P9 => unnamed_net34,
      P10 => unnamed_net17,
      P8 => unnamed_net35,
      
      P4 => unnamed_net36,
      P5 => unnamed_net17,
      P6 => unnamed_net37,
      
      P1 => unnamed_net38,
      P2 => unnamed_net17,
      P3 => unnamed_net39,
      
      P12 => Vcc,
      P13 => unnamed_net17,
      P11 => unnamed_net41,
      P14 => Vcc,
      P7 => GND);

  U10 : hc7486
    PORT MAP (
      P1 => unnamed_net11,
      P2 => unnamed_net15,
      P3 => unnamed_net32,
      
      P4 => unnamed_net13,
      P5 => unnamed_net15,
      P6 => unnamed_net33,
      
      P9 => unnamed_net22,
      P10 => Vcc,
      P8 => unnamed_net55,
      
      P12 => Vcc,
      P13 => unnamed_net53,
      P11 => unnamed_net54,
      P14 => Vcc,
      P7 => GND);

  U9 : hc7486
    PORT MAP (
      P1 => unnamed_net1,
      P2 => unnamed_net15,
      P3 => unnamed_net28,
      
      P4 => unnamed_net3,
      P5 => unnamed_net15,
      P6 => unnamed_net29,
      
      P9 => unnamed_net5,
      P10 => unnamed_net15,
      P8 => unnamed_net30,
      
      P12 => unnamed_net7,
      P13 => unnamed_net15,
      P11 => unnamed_net31,
      P14 => Vcc,
      P7 => GND);

  U1 : hc74163
    PORT MAP (
      P3 => GND,
      P14 => unnamed_net22,
      P4 => GND,
      P13 => unnamed_net23,
      P5 => GND,
      P12 => unnamed_net24,
      P6 => GND,
      P11 => unnamed_net25,
      P7 => Vcc,
      P15 => unnamed_net26,
      P10 => Vcc,
      P2 => unnamed_net27,
      P1 => Vcc,
      P9 => Vcc,
      P16 => Vcc,
      P8 => GND);

  U6 : hc74273
    PORT MAP (
      P11 => unnamed_net21,
      P3 => unnamed_net2,
      P4 => unnamed_net4,
      P7 => unnamed_net6,
      P8 => unnamed_net8,
      P13 => unnamed_net12,
      P14 => unnamed_net14,
      P17 => unnamed_net16,
      P18 => unnamed_net18,
      P1 => Vcc,
      P2 => unnamed_net1,
      P5 => unnamed_net3,
      P6 => unnamed_net5,
      P9 => unnamed_net7,
      P12 => unnamed_net11,
      P15 => unnamed_net13,
      P16 => unnamed_net15,
      P19 => unnamed_net17,
      P20 => Vcc,
      P10 => GND);

  U4 : hc74283
    PORT MAP (
      P5 => unnamed_net11,
      P4 => unnamed_net12,
      P3 => unnamed_net13,
      P1 => unnamed_net14,
      P14 => unnamed_net15,
      P13 => unnamed_net16,
      P12 => unnamed_net17,
      P10 => unnamed_net18,
      P6 => unnamed_net9,
      P9 => unnamed_net19,
      P2 => GND,
      P15 => unnamed_net20,
      P11 => GND,
      P7 => unnamed_net10,
      P16 => Vcc,
      P8 => GND);

  U5 : hc74283
    PORT MAP (
      P5 => unnamed_net1,
      P4 => unnamed_net2,
      P3 => unnamed_net3,
      P1 => unnamed_net4,
      P14 => unnamed_net5,
      P13 => unnamed_net6,
      P12 => unnamed_net7,
      P10 => unnamed_net8,
      P6 => unnamed_net9,
      P9 => unnamed_net10,
      P2 => GND,
      P15 => unnamed_net9,
      P11 => GND,
      P7 => GND,
      P16 => Vcc,
      P8 => GND);

  vcc <= '1';
  gnd <= '0';

  

-- Signal assignment part
END netlist;
